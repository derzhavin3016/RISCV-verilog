`include "consts.v"

module datapath (input clk, reset,
                     input memtoreg, pcsrc,
                     input [1:0] alusrc,
                     input regwrite, jump,
                     input [3:0] alucontrol,
                     output zero,
                     output [31:0] pc,
                     input [31:0] instr,
                     output [31:0] aluout, writedata,
                     input [31:0] readdata
                    );
    wire [4:0] writereg;
    wire [31:0] pcnext, pcnextbr, pcplus4, pcbranch;
    wire [31:0] imm;
    wire [31:0] srca, srcb;
    wire [31:0] result;
    // next PC logic
    flopr #(32) pcreg(clk, reset, pcnext, pc);
    adder pcadd1(pc, 32'd4, pcplus4);
    adder pcadd2(pcplus4, immsh, pcbranch);

    mux2 #(32) pcbrmux(pcplus4, pcbranch, pcsrc, pcnextbr);
    mux2 #(32) pcmux(pcnextbr, {pcplus4[31:28], instr[25:0], 2'b00}, jump, pcnext);

    // register file logic
    immSel immsel(instr, imm);
    regfile rf(clk, regwrite, instr[25:21],
               instr[20:16], writereg,
               result, srca, writedata);
    mux2 #(5) wrmux(instr[20:16], instr[15:11], regdst, writereg);
    mux2 #(32) resmux(aluout, readdata, memtoreg, result);
    signext se(instr[15:0], imm);

    // ALU logic
    mux4 #(32) srcbmux(writedata, imm, alusrc, srcb);
    alu alu(srca, srcb, alucontrol, aluout, zero);
endmodule
